library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ram_tempos is
   port (       
       clk          : in  std_logic;
       endereco     : in  std_logic_vector(7 downto 0);
       dado_entrada : in  std_logic_vector(13 downto 0);--tempo de reacao do jogador
       we           : in  std_logic;
       ce           : in  std_logic;
       dado_saida   : out std_logic_vector(13 downto 0)
    );
end entity ram_tempos;

architecture ram_mif of ram_tempos is
  type   arranjo_memoria is array(0 to 255) of std_logic_vector(13 downto 0);
  signal memoria : arranjo_memoria;
  
  -- Configuracao do Arquivo MIF
  attribute ram_init_file: string;
  attribute ram_init_file of memoria: signal is "ram_tempos_inicial.mif";
  
begin

  process(clk)
  begin
    if (clk = '1' and clk'event) then
          if ce = '0' then -- dado armazenado na subida de "we" com "ce=0"
           
              -- Detecta ativacao de we (ativo baixo)
              if (we = '0') 
                  then memoria(to_integer(unsigned(endereco))) <= dado_entrada;
              end if;
            
          end if;
      end if;
  end process;

  -- saida da memoria
  dado_saida <= memoria(to_integer(unsigned(endereco)));
  
end architecture ram_mif;

-- Dados iniciais (para simulacao com Modelsim) 
architecture ram_modelsim of ram_tempos is
  type   arranjo_memoria is array(0 to 255) of std_logic_vector(13 downto 0);
  signal memoria : arranjo_memoria := ( "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
													 "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000",
                                        "00000000000000");
  
begin

  process(clk)
  begin
    if (clk = '1' and clk'event) then
          if ce = '0' then -- dado armazenado na subida de "we" com "ce=0"
              -- Detecta ativacao de we (ativo baixo)
              if (we = '0') 
                  then memoria(to_integer(unsigned(endereco))) <= dado_entrada;
              end if;
            
          end if;
      end if;
  end process;

  -- saida da memoria
  dado_saida <= memoria(to_integer(unsigned(endereco)));

end architecture ram_modelsim;